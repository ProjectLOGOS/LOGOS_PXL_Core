From Coq Require Import Program.

(* TODO: Restore full imports once module path resolution is fixed *)
(* From PXLs Require Import PXLv3. *)
(* Require Import modules.chronopraxis.substrate.ChronoAxioms *)
(*                modules.chronopraxis.theorems.MetaTheorems. *)

(* Standalone definitions for compilation *)
Inductive form : Type :=
| Bot : form
| Atom : nat -> form
| Impl : form -> form -> form
| Conj : form -> form -> form
| Disj : form -> form -> form
| Neg : form -> form
| Box : form -> form
| Dia : form -> form.

Parameter Gamma : Type.
Definition can_world := {gamma : Gamma | True}.
Parameter forces : can_world -> form -> Prop.
Parameter In_set : Gamma -> form -> Prop.

Set Implicit Arguments.

(* Syntactic predicate: no Box/Dia inside φ *)
Fixpoint modal_free (φ: form) : Prop :=
  match φ with
  | Bot | Atom _ => True
  | Impl a b | Conj a b | Disj a b => modal_free a /\ modal_free b
  | Neg a => modal_free a
  | Box _ | Dia _ => False
  end.

(* Truth lemma bridge - would use kernel's truth lemma when available *)
Parameter truth_lemma : forall (w: can_world) (φ: form), 
  forces w φ <-> In_set (proj1_sig w) φ.

(* Semantic collapse: for modal-free φ, forces ignores R and matches base truth in Γ. *)
Lemma forces_modal_free_eq_membership :
  forall (w: can_world) (φ: form),
    modal_free φ ->
    (forces w φ <-> In_set (proj1_sig w) φ).
Proof.
  (* By your constructive Truth Lemma, forces w φ <-> In_set Γ φ for all φ.
     This lemma is stated to expose explicitly the modal_free precondition used later. *)
  intros w φ _. apply truth_lemma.
Qed.
