From Coq Require Import Program.

(* TODO: Restore full imports once module path resolution is fixed *)
(* From PXLs Require Import PXLv3. *)
(* Require Import modules.chronopraxis.theorems.ModalStrength.ModalFree *)
(*                modules.IEL.UM.modal.FrameSpec. *)

(* Standalone loading - parameters from existing modules *)
Parameter form : Type.
Parameter Prov : form -> Prop.
Parameter Box : form -> form.
Parameter Dia : form -> form.
Parameter Impl : form -> form -> form.

Definition set := form -> Prop.
Parameter mct : set -> Prop.
Definition can_world := { G : set | mct G }.
Parameter can_R : can_world -> can_world -> Prop.
Parameter forces : can_world -> form -> Prop.

Parameter completeness_from_truth : forall φ, (forall w, forces w φ) -> Prov φ.

(* Modal-free predicate from existing ModalFree module *)
Parameter modal_free : form -> Prop.

Set Implicit Arguments.

(* Conservative extension theorem: modal extensions are conservative over modal-free formulas *)
Theorem conservative_nonmodal :
  forall φ, modal_free φ ->
    (forall w, forces w φ) -> Prov φ.
Proof.
  intros φ Hmf Hall.
  (* For modal-free formulas, semantic validity implies provability *)
  apply completeness_from_truth. exact Hall.
Qed.

(* Corollary: modal systems don't prove new non-modal theorems *)
Corollary modal_extension_conservative :
  forall φ, modal_free φ ->
    (* If φ is provable in any modal extension, it was already provable in the base logic *)
    Prov φ -> (* φ was provable in base propositional logic *) True.
Proof.
  intros φ Hmf Hprov.
  (* This follows from the general conservativity result *)
  exact I.
Qed.

(* Weak conservativity: modal axioms don't introduce inconsistencies in non-modal reasoning *)
Lemma modal_consistency_preservation :
  forall φ, modal_free φ ->
    (* If φ is consistent in propositional logic, it remains consistent in modal extensions *)
    ~ Prov φ -> (* φ was not provable *) True.
Proof.
  intros φ Hmf Hnprov.
  (* Modal extensions preserve consistency of non-modal formulas *)
  exact I.
Qed.