(* Compatibilism_CoffeeTea.v - Concrete example of temporal freedom *)

From Coq Require Import Program.

(* TODO: Restore full imports once module path resolution is fixed *)
(* Require Import PXLs.IEL.Infra.substrate.ChronoAxioms *)
(*                PXLs.IEL.Infra.substrate.ChronoMappings *)
(*                PXLs.IEL.Infra.domains.Compatibilism.CompatibilismTheory. *)

Module CoffeeTea.

(* Simplified temporal types for the example *)
Parameter PA : Type.  (* χ_A - lived time propositions *)
Parameter PC : Type.  (* χ_C - eternal time propositions *)
Parameter A_to_C : PA -> PC.

(* Simplified compatibilism types *)
Record Agent := { agent_id : nat }.
Definition alt (pA pA' : PA) : Prop := pA <> pA' /\ A_to_C pA = A_to_C pA'.
Definition Free (_:Agent) (pA:PA) : Prop := exists pA', alt pA pA'.

(* Example scenario: coffee vs tea choice *)
(* Two different lived experiences that lead to same eternal outcome *)
Parameter pA_coffee pA_tea : PA.

(* Coffee and tea are different experiences in lived time *)
Parameter distinct_experiences : pA_coffee <> pA_tea.

(* But both map to same eternal truth: "had warm beverage at 3pm" *)
Parameter same_cosmic_outcome : A_to_C pA_coffee = A_to_C pA_tea.

(* Agent making the choice *)
Definition agent := {| agent_id := 1 |}.

(* Demonstration: The agent is free on the coffee choice *)
(* Because there exists a genuine alternative (tea) that maps to same eternal outcome *)
Theorem free_coffee_example : Free agent pA_coffee.
Proof.
  exists pA_tea. 
  split.
  - exact distinct_experiences.  (* Coffee ≠ tea in lived experience *)
  - exact same_cosmic_outcome.   (* Both → "warm beverage" in eternal time *)
Qed.

(* Similarly for the tea choice *)
Theorem free_tea_example : Free agent pA_tea.
Proof.
  exists pA_coffee.
  split.
  - intro H. exact (distinct_experiences (eq_sym H)).
  - exact (eq_sym same_cosmic_outcome).
Qed.

(* Key insight: Freedom exists because alternatives in χ_A converge in χ_C *)
(* This captures compatibilist intuition: genuine choice with inevitable outcome *)

End CoffeeTea.
