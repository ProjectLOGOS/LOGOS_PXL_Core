From Coq Require Import Program.

(* TODO: Restore full imports once module path resolution is fixed *)
(* From PXLs Require Import PXLv3. *)
(* Require Import PXLs.IEL.Infra.theorems.ModalStrength.S4Overlay *)
(*                PXLs.IEL.Infra.theorems.ModalStrength.S5Overlay *)
(*                PXLs.IEL.Infra.theorems.ModalStrength.ModalAxiomsSound. *)

(* Standalone loading for compilation - using direct compilation approach *)
Parameter form : Type.
Parameter Prov : form -> Prop.
Parameter Box : form -> form.
Parameter Dia : form -> form.
Parameter Impl : form -> form -> form.

(* Parameters for the proven theorems *)
Parameter provable_T : forall φ, Prov (Impl (Box φ) φ).
Parameter provable_4 : forall φ, Prov (Impl (Box φ) (Box (Box φ))).
Parameter provable_5 : forall φ, Prov (Impl (Dia φ) (Box (Dia φ))).
Parameter provable_B : forall φ, Prov (Impl φ (Box (Dia φ))).

Goal True. exact I. Qed.

(* Verify that all modal axiom schemata are available *)
Check provable_T.     (* T axiom: □φ → φ *)
Check provable_4.     (* 4 axiom: □φ → □□φ *)
Check provable_5.     (* 5 axiom: ◇φ → □◇φ *)
Check provable_B.     (* B axiom: φ → □◇φ *)

(* Example: instantiate the axioms with a concrete formula *)
Parameter A : nat.
Parameter Atom : nat -> form.
Definition example_atom := Atom A.

(* The axioms apply to any formula, including our example *)
Example T_instance : Prov (Impl (Box example_atom) example_atom).
Proof. apply provable_T. Qed.

Example four_instance : Prov (Impl (Box example_atom) (Box (Box example_atom))).
Proof. apply provable_4. Qed.

Example five_instance : Prov (Impl (Dia example_atom) (Box (Dia example_atom))).
Proof. apply provable_5. Qed.

Example B_instance : Prov (Impl example_atom (Box (Dia example_atom))).
Proof. apply provable_B. Qed.

(* Demonstrate that we have the complete S4 and S5 axiomatizations *)
Lemma S4_axioms_complete : forall φ, 
  Prov (Impl (Box φ) φ) /\                    (* T *)
  Prov (Impl (Box φ) (Box (Box φ))).          (* 4 *)
Proof.
  intro φ. split.
  - apply provable_T.
  - apply provable_4.
Qed.

Lemma S5_axioms_complete : forall φ,
  Prov (Impl (Box φ) φ) /\                    (* T *)
  Prov (Impl (Box φ) (Box (Box φ))) /\        (* 4 *)
  Prov (Impl (Dia φ) (Box (Dia φ))).          (* 5 *)
Proof.
  intro φ. split; [| split].
  - apply provable_T.
  - apply provable_4.
  - apply provable_5.
Qed.

(* Alternative S5 axiomatization using Brouwer axiom *)
Lemma S5_Brouwer_axioms : forall φ,
  Prov (Impl (Box φ) φ) /\                    (* T *)
  Prov (Impl φ (Box (Dia φ))).                (* B - Brouwer axiom *)
Proof.
  intro φ. split.
  - apply provable_T.
  - apply provable_B.
Qed.
